module coder83(I,O)
{
    input
}