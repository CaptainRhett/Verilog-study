module basic_rs_latch(R,S,Q,NQ);
    input R;
    input S;
    wire Q;
    wire NQ;
    
