module code_88_logic;
    input [7:0]i;
    output [2:0]o;