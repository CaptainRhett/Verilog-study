module adder(A,B,Y);
    input [3:0]A;
    input [3:0]B;
    output [3:0]Y;
    wire [3:0]Y;
    assing Y = A + B;
endmodule: